-- hps.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity hps is
	port (
		h2f_loan_io_in                   : out   std_logic_vector(66 downto 0);                    -- h2f_loan_io.in
		h2f_loan_io_out                  : in    std_logic_vector(66 downto 0) := (others => '0'); --            .out
		h2f_loan_io_oe                   : in    std_logic_vector(66 downto 0) := (others => '0'); --            .oe
		hps_io_hps_io_gpio_inst_LOANIO49 : inout std_logic                     := '0';             --      hps_io.hps_io_gpio_inst_LOANIO49
		hps_io_hps_io_gpio_inst_LOANIO50 : inout std_logic                     := '0';             --            .hps_io_gpio_inst_LOANIO50
		hps_io_hps_io_gpio_inst_LOANIO53 : inout std_logic                     := '0';             --            .hps_io_gpio_inst_LOANIO53
		hps_io_hps_io_gpio_inst_LOANIO54 : inout std_logic                     := '0';             --            .hps_io_gpio_inst_LOANIO54
		memory_mem_a                     : out   std_logic_vector(14 downto 0);                    --      memory.mem_a
		memory_mem_ba                    : out   std_logic_vector(2 downto 0);                     --            .mem_ba
		memory_mem_ck                    : out   std_logic;                                        --            .mem_ck
		memory_mem_ck_n                  : out   std_logic;                                        --            .mem_ck_n
		memory_mem_cke                   : out   std_logic;                                        --            .mem_cke
		memory_mem_cs_n                  : out   std_logic;                                        --            .mem_cs_n
		memory_mem_ras_n                 : out   std_logic;                                        --            .mem_ras_n
		memory_mem_cas_n                 : out   std_logic;                                        --            .mem_cas_n
		memory_mem_we_n                  : out   std_logic;                                        --            .mem_we_n
		memory_mem_reset_n               : out   std_logic;                                        --            .mem_reset_n
		memory_mem_dq                    : inout std_logic_vector(39 downto 0) := (others => '0'); --            .mem_dq
		memory_mem_dqs                   : inout std_logic_vector(4 downto 0)  := (others => '0'); --            .mem_dqs
		memory_mem_dqs_n                 : inout std_logic_vector(4 downto 0)  := (others => '0'); --            .mem_dqs_n
		memory_mem_odt                   : out   std_logic;                                        --            .mem_odt
		memory_mem_dm                    : out   std_logic_vector(4 downto 0);                     --            .mem_dm
		memory_oct_rzqin                 : in    std_logic                     := '0'              --            .oct_rzqin
	);
end entity hps;

architecture rtl of hps is
	component hps_hps is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_loan_in               : out   std_logic_vector(66 downto 0);                    -- in
			h2f_loan_out              : in    std_logic_vector(66 downto 0) := (others => 'X'); -- out
			h2f_loan_oe               : in    std_logic_vector(66 downto 0) := (others => 'X'); -- oe
			mem_a                     : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                    : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                    : out   std_logic;                                        -- mem_ck
			mem_ck_n                  : out   std_logic;                                        -- mem_ck_n
			mem_cke                   : out   std_logic;                                        -- mem_cke
			mem_cs_n                  : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                 : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                 : out   std_logic;                                        -- mem_cas_n
			mem_we_n                  : out   std_logic;                                        -- mem_we_n
			mem_reset_n               : out   std_logic;                                        -- mem_reset_n
			mem_dq                    : inout std_logic_vector(39 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                   : inout std_logic_vector(4 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                 : inout std_logic_vector(4 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                   : out   std_logic;                                        -- mem_odt
			mem_dm                    : out   std_logic_vector(4 downto 0);                     -- mem_dm
			oct_rzqin                 : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_gpio_inst_LOANIO49 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO49
			hps_io_gpio_inst_LOANIO50 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO50
			hps_io_gpio_inst_LOANIO53 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO53
			hps_io_gpio_inst_LOANIO54 : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO54
			h2f_rst_n                 : out   std_logic                                         -- reset_n
		);
	end component hps_hps;

begin

	hps : component hps_hps
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			h2f_loan_in               => h2f_loan_io_in,                   -- h2f_loan_io.in
			h2f_loan_out              => h2f_loan_io_out,                  --            .out
			h2f_loan_oe               => h2f_loan_io_oe,                   --            .oe
			mem_a                     => memory_mem_a,                     --      memory.mem_a
			mem_ba                    => memory_mem_ba,                    --            .mem_ba
			mem_ck                    => memory_mem_ck,                    --            .mem_ck
			mem_ck_n                  => memory_mem_ck_n,                  --            .mem_ck_n
			mem_cke                   => memory_mem_cke,                   --            .mem_cke
			mem_cs_n                  => memory_mem_cs_n,                  --            .mem_cs_n
			mem_ras_n                 => memory_mem_ras_n,                 --            .mem_ras_n
			mem_cas_n                 => memory_mem_cas_n,                 --            .mem_cas_n
			mem_we_n                  => memory_mem_we_n,                  --            .mem_we_n
			mem_reset_n               => memory_mem_reset_n,               --            .mem_reset_n
			mem_dq                    => memory_mem_dq,                    --            .mem_dq
			mem_dqs                   => memory_mem_dqs,                   --            .mem_dqs
			mem_dqs_n                 => memory_mem_dqs_n,                 --            .mem_dqs_n
			mem_odt                   => memory_mem_odt,                   --            .mem_odt
			mem_dm                    => memory_mem_dm,                    --            .mem_dm
			oct_rzqin                 => memory_oct_rzqin,                 --            .oct_rzqin
			hps_io_gpio_inst_LOANIO49 => hps_io_hps_io_gpio_inst_LOANIO49, --      hps_io.hps_io_gpio_inst_LOANIO49
			hps_io_gpio_inst_LOANIO50 => hps_io_hps_io_gpio_inst_LOANIO50, --            .hps_io_gpio_inst_LOANIO50
			hps_io_gpio_inst_LOANIO53 => hps_io_hps_io_gpio_inst_LOANIO53, --            .hps_io_gpio_inst_LOANIO53
			hps_io_gpio_inst_LOANIO54 => hps_io_hps_io_gpio_inst_LOANIO54, --            .hps_io_gpio_inst_LOANIO54
			h2f_rst_n                 => open                              --   h2f_reset.reset_n
		);

end architecture rtl; -- of hps
